sngl single                                                                                         L1-1        `�Q@L2-2        5~�@L1-1-END    ��N@L2-2-END    H��@
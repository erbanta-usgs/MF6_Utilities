cont double  40                                                                                        RIV1-3-1                                RIV1-4-2                                RIV1-5-3                                RIV1-5-4                                RIV2-7-4                                RIV2-7-5                                RIV2-9-6                                      �?����:�@@��Po�@ ۸C}��@�k�E��@ ��n>��@���i��@�i8���BFUUUUUU�?�\�U+�@�]�i�ơ@ �-vZ�@��ud��@P���r�@ K���@�i8���BF�������?��:�v�@@���7�@���XK��@P��؍٣@�����@�z=��@�i8���BF�������?�Y�"��@��Dt,]�@��̓�@�i�*%�@p�K��@���h��@�i8���BFTUUUUU�?@�u7�@�w�O���@�s��O<�@ �F�:p�@�5�Rvߡ@���쾈�@�i8���BF�������?�FҿT�@p�qr�@����@��*���@P��e�ݡ@�ʓ���@�i8���BF�������?�g�1���@з�5�:�@@:�i"Ц@@E2R��@��8'ܡ@�=��j��@�i8���BFSUUUUU�? ���/�@І|���@0!�K:�@P�� N�@�K�v�ڡ@���@�i8���BF�������? �hh.�@�B��˪@o�Y�a�@@j����@� Q��ء@ ׼���@�i8���BF�������?�ӵuu�@0]Bz�@��M�ɩ�@��ԃS߬@�J�K;ס@ *�x��@�i8���BFRUUUUU�?��I��@0�^R�Z�@0�u1B�@ 2�'�@�(��ա@�P��~�@�i8���BF�������?���f��@�:�C��@К�!08�@`�ݥ]n�@�R��ӡ@@���-}�@�i8���BF�������?Pp�TH�@Ѕ�Y�@�ۨ�~�@�M�D�Z�@�X7WXҡ@����{�@�i8���BF������ @ ��h�F�@�7�s��@P��~nį@�u���@�����@ Ʉh4e�@�i8���BFTUUUUU@PFM�@h���8�@@�z���@pϮ"p��@�t�o·�@PܶO�a�@�i8���BF������@��d*2��@�8*6۱@����D'�@о�-�B�@�I��{��@P7瓖^�@�i8���BF������@��.-�@�ae�1}�@��z7eɱ@0���E�@�)��6��@��I�I[�@�i8���BFUUUUUU@����β@h�N���@0S�Ak�@(-IJ��@�é�@�Z���W�@�i8���BF      @pDF�o�@��x�^��@��_J��@��y
)�@P[�3���@`�,��T�@�i8���BF������@P�����@0I�X�a�@h�G@/��@����ʴ@�:N�r��@��\KfQ�@�i8���BFVUUUUU@��鞱�@�;X/�@��Z�@O�@�8�k�@ k��6��@0G�	N�@�i8���BF     @��2R�@��j+��@X�|�@�h��@������@@w
#�J�@�i8���BF������@ �J�Z�@�>�6�C�@E����@�>�bi��@0s�ŝ�@0�ߕG�@�i8���BFWUUUUU@8K�T��@xД���@`�x��0�@�Ù��M�@Ъ�����@0yYQD�@�i8���BF     @�n�2�@ض�����@�fX�ж@X��X�@="[��@�H��A�@�i8���BF������@^D�T�@�K�:��@؍rށ�@HF�y��@���׫@p�uh��@�i8���BFXUUUUU	@�v��(��@�z.�K�@�J �☶@ ��W쵷@��)Sҫ@��J=)}�@�i8���BF     
@h&	�㟶@hh�wf�@h"�hl>�@@���\[�@�˿Y,̫@`�u)>w�@�i8���BF������
@�y�v�E�@8�h9��@�9>>�@H���� �@@�cXƫ@��O�Uq�@�i8���BFYUUUUU@��O��@�PP�4=�@���)���@���Ӷ��@��/ׇ��@���#ok�@�i8���BF     @�����@ td�X�@hS���/�@(K��L�@��E����@@�F�e�@�i8���BF������@ /%k^8�@X������@����#ִ@`2�H��@`"��@�����_�@�i8���BFZUUUUU@��F}�޴@�v��0�@��Mu|�@�P�(阵@���+��@��%��Y�@�i8���BF     @8$&���@�+��ִ@H?���"�@XQ�1J?�@���Fk��@P�[�S�@�i8���BF������@��gO[,�@@zy}�@ L�ɳ@�ϑ	��@�ƾ���@�x�qN�@�i8���BF[UUUUU@�>�Sӳ@��,e$�@P��Xp�@x�Y7���@0H����@ڜPIH�@�i8���BF     @(x��sz�@"E�x˳@ ��H�@H�NxZ3�@��G?��@ ��vB�@�i8���BFXUUUUU@�hv>�6�@þ�@`��?<Ӳ@��ҝ:�@PN	yz#�@@�z��ͯ@�i8���BF������@��sє�@@�%˒X�@����*��@�QY���@P1�� �@0��X�ǯ@�i8���BF     @X�֣�ز@(�8L�)�@�}�;.u�@H����@�p
k��@�6G���@�i8���BFWUUUUU@���婲@�;�g���@���UGF�@`�[�b�@�>��z�@���Q���@�i8���BF������@`���-{�@��_,̲@�j��u�@��&=3�@�7�.
�@�;6��@�i8���BF     @���L�@؇����@�P� ��@����r�@�����@P�;̭�@�i8���BFVUUUUU@���\��@���R�n�@ w�a��@ .�ղ@�X�����@�A�me��@�i8���BF������@��L���@��4�@�@f8�~��@Шu���@�Y��^��@`&���@�i8���BF      @X�� ��@@�!�#�@@��]�@ E�5�x�@��r�"�@�������@�i8���BFUUUUUU@�Ø�ђ�@��
��@�}2A�.�@ F6�J�@@Xu���@@�SN��@�i8���BF������@HQɠ�d�@���U���@8���E �@��&ػ�@@����@p������@�i8���BF������@�oBr6�@ `�|��@�Ǿ:Ұ@�#P�o�@0��ެ@@@Ii���@�i8���BFTUUUUU@Z�a�@�[Y�nY�@pI0ݣ�@ȝ�7��@���8[ج@�׻�Q��@�i8���BF������@�B�meڰ@�!v+�@(���u�@8����@��W�2Ҭ@��d�{�@�i8���BF������@�/�}��@8�����@@�=�G�@�
e�c�@�G)�̬@p{�j�t�@�i8���BFSUUUUU@0/��~�@�bh��ϰ@x�c��@p�$�5�@��Gf�Ŭ@�_�wn�@�i8���BF������@��wm�P�@�����@0K�<د@H�P)�@ ֱ�ӿ�@ ��5h�@�i8���BF������@X�]B#�@8/�bt�@��W��|�@����Xٰ@���⻹�@P0n�a�@�i8���BFRUUUUU@�a�JY�@����F�@P��~%!�@�វ��@���p���@0���[�@�i8���BF������@�5/pV��@ �TU�@�e D�Ů@H"w�}�@PU�3���@@����U�@�i8���BF������@`h$|5�@0���ׯ@����j�@�UNbP�@@�뮋��@�+AOO�@�i8���BFQUUUUU@ ��\�ڮ@��3}�@p�F��@�f�'�"�@�.z��@P�L� I�@�i8���BF������@�,S�@��@��ı�"�@0��I��@ �?}��@ 89����@���o�B�@�i8���BF������@@����%�@�[GG`Ȯ@��S`�Z�@�KokH��@�6�����@�����<�@�i8���BFPUUUUU@04��٭@ z��|�@��'7�@0��˯C�@ ���W�@��ʖN��@�i8���BF������@p�;3��@�1���=�@@l��Ϭ@`�'%�@~"K�Q�@�+�|���@�i8���BF������@ �ٔ�\�@ 2)���@�+9Oe��@��@�Ʈ@�1��dK�@��a�@�i8���BFOUUUUU@�G���@�������@`o\'S�@��/f��@����E�@�Zǅ��@�i8���BF������@pH�i��@Pi�?���@p�Z��@�Ȁ1J�@P�>�@�B�ކ�@�i8���BF������@�紹���@�ٟ��E�@�H��֫@p����@�|���8�@���߯@�i8���BFNUUUUU@�g�/e�@ �|B;�@P���@���έ@��czh2�@0t-�د@�i8���BF������@��G��'�@��ͣʬ@ ��ME[�@ Lr�7��@���3,�@\�Uү@�i8���BF������@ �p���@�*e(��@ 0z��@0ʇ�qR�@�X&�@��vN�˯@�i8���BFMUUUUU@��{��@���O�@�,Y��ߪ@ S{���@�67n��@0�F��ů@�i8���BF������@�^�� o�@ #���@�Q�À��@��A;׬@ ����@���L��@�i8���BF������@���1�@�r$^ի@`��>!e�@���ș�@@�;���@@}����@�i8���BFLUUUUU@��s���@�noR��@`����'�@��BPq\�@p���i�@pi����@�i8���BF������@�Ҵ-���@���a[�@�~	���@e^�4�@PC�UL�@ ��^��@�i8���BF������@��;�z�@��(k��@Pi�ץ��@ ���@�Z�r3�@�$�Y��@�i8���BFKUUUUU@��&'�=�@��\���@p_L��p�@��(B��@`�V-��@��=՟�@�i8���BF������@�3�^@�@ 9��4��@�Qږ�3�@P��%h�@���#��@P�����@�i8���BF������@ ���ĩ@���αh�@迳 ��@0j�YW+�@`Y��@�ѥ6[��@�i8���BFJUUUUU@�� �#��@�e�J,�@0����@W�J��@����@���!��@�i8���BF������@��ƽK�@�v�N��@�)\�}�@���
��@�v>d��@ࣵ�솯@�i8���BF������@���r�@�<��˳�@�Rl#�A�@��IG�u�@@���ܬ@>fX���@�i8���BFIUUUUU@0�BӨ@0���w�@@�>�@ 4$%*9�@��5l�֬@�Tv�z�@�i8���BF������@�-m,��@PS6u�;�@ �^	ɧ@0Zd0���@��ߖ�Ь@P���jt�@�i8���BF������@P-gj1[�@��3����@k��@О�����@�A�Jˬ@@� Fn�@�i8���BF�����* @ B�P�@�'��Ĩ@@�[��P�@0`�ࣄ�@pmSŬ@0wq#h�@�i8���BFOUUUUU @�:Ċ�@���g��@��W��@0>A�H�@�_S,��@���b�@�i8���BF����� @`���ާ�@ d���L�@`��=٦@���U��@`Kf�B��@���I�[�@�i8���BF������ @�РjMl�@�3o_�@ 0�����@@/�y
Ѩ@ p�V]��@`�׺�U�@�i8���BFPUUUU� @���1�0�@��?d֧@�,r��a�@�p�gb��@ o�X|��@P�e�O�@�i8���BF������ @��1y��@��O����@P��{&�@ ��r�Y�@�KZ����@`�sܳI�@�i8���BF�����*!@ ��G6��@��IA�_�@�9*�@`��&`�@�g�ġ�@�ݪ�C�@�i8���BFQUUUUU!@P��X�@p�ی$�@@Б@ѯ�@`Փ��@�hYG@�B�͞=�@�i8���BF�����!@@S�X�C�@��∙�@��s�t�@��c�ŧ�@pjh���@�Er̚7�@�i8���BF������!@���J		�@@(Z���@��8��9�@`��a�l�@�y�M��@�e:�1�@�i8���BFRUUUU�!@0�,.Υ@�^Kt�@�D�����@0�f��1�@`pF���@P���+�@�i8���BF������!@��l��@0c�5\9�@@�oi�ä@�QL����@���Q���@P,���%�@�i8���BF�����*"@@�*�J�@pz
#��@P�f`	{�@`��୦@��0��@�a*���@�i8���BFSUUUUU"@����@p:xѶ��@���c�$�@��H�PW�@ QY	Q �@�:�s��@�i8���BF�����"@@i�t��@p��٦D�@�=�@Σ@�c�� �@�0����@0֕�ۛ�@�i8���BF������"@����tH�@��@��@`G��x�@��&����@������@@;�G��@�i8���BFTUUUU�"@ �Vș�@�#_����@ �7;"�@ Ʋ��T�@ ?Hi$��@�rh����@�i8���BF������"@p��%䜣@ �u�VC�@ଁ-̢@��5����@ ����@��X�%��@�i8���BF�����*#@�&�|SG�@�����@P1��pv�@�2�岨�@@�]Sg�@�
�o���@�i8���BFUUUUUU#@��D���@p�����@0�ZM� �@ ��fS�@0TD�@�p ���@�i8���BF     �#@PUˇ���@0ݕ0TC�@�3�fˡ@X�v��@�^�v��@��}��@�i8���BF������#@`��~G�@�UU}G�@���'v�@���+��@0{�~Z�@ �����@�i8���BFVUUUU�#@��_��@ЎE�_��@�`�� �@P9���R�@ ѱZ�@ �w5s�@�i8���BF     $@`ó9���@���A�D�@��X�ˠ@@��=���@P�h�ަ@���G�{�@�i8���BF�����*$@�݁�H�@��U��@P]Եw�@�G����@��%�cۦ@�-�ox�@�i8���BFWUUUUU$@���b��@�ȏ���@�{UR"�@� F��S�@p;e�ئ@�)�t�@�i8���BF    �$@�π����@��o�+G�@����v��@ �:��@P�;��Ԧ@L��pq�@�i8���BF������$@@Tvb�K�@�_X(��@ �`T��@��2���@0�;}Ѧ@}��m�@�i8���BFXUUUU�$@ ��D�@ "U�Ꞡ@`���I�@���IV�@���,5Φ@0&b�~j�@�i8���BF     %@ Q�G�@��Q��J�@�9�]���@�vG�@@���ʦ@ �d	g�@�i8���BF�����*%@ �$�X��@�_��q�@ �%Г��@�hO魠@@�Ä�Ǧ@�+��c�@�i8���BFYUUUUU%@� Do���@�%N+G�@�X-�Q�@Զ9�Y�@���iĦ@��~�!`�@�i8���BF    �%@��>%�P�@�G��+��@�>�zP��@�,"�@�6�(��@��7 �\�@�i8���BF������%@ ٜ�٩�@����r��@�IR*�@�l���d�@0�û꽦@�a�?DY�@�i8���BFZUUUU�%@�X��=�@`]wS�@�}��+\�@`ri���@�s�����@`��U�@�i8���BF     &@��>��\�@�,�֬�@ �wĄ��@������@ }�w��@���4tR�@�i8���BF�����*&@�x ��@ ᙉR�@`��HZ�@ ���z��@ �ŕ"P�@�i�AA�@�i8���BF[UUUUU&@@6����@�E�ScB�@@y�SJ�@@��Vv��@��/	�O�@@a{S�@�@�i8���BF    �&@���-��@���)�2�@`�߯j:�@ R }��@ x�$[O�@@�}�U@�@�i8���BF������&@ ?���њ@@,�D#�@@֖��*�@�2�����@ ���N�@ ")�?�@�i8���BF\UUUU�&@�E�E@`�����@�����@`ɯ�{�@���B�N�@���?�@�i8���BF     '@@5RD��@ fc�H�@���
�@�^^|�k�@ {��CN�@`JӀI?�@�i8���BF�����*'@�\Q�t��@��g����@`��$��@@`P��[�@�e���M�@�b���>�@�i8���BF]UUUUU'@`�6���@@���k�@�a0f�@`1L�@`.���M�@ �U�>�@�i8���BF    �'@�U�z삚@���\֛@`B� �ۘ@`�q;k<�@ �i�5M�@�#[A>�@�i8���BF������'@��e�2s�@@�o��ƛ@ X�>�˘@ �J�,�@ ��<�L�@0�.�=�@�i8���BF^UUUU�'@`�oR�c�@@��R��@@�G�V��@ �P���@@����L�@�=��=�@�i8���BF	     (@����S�@��8��@������@`%��I�@@��1L�@ �c�C=�@�i8���BF�����*(@� 9�/D�@�wD���@ �F@��@�Q���@��S�K�@ c���<�@�i8���BF_UUUUU(@ �%��4�@�rt��@ %ⴆ��@ \�A��@@K�W�K�@P��X�<�@�i8���BF
    �(@@8��$�@���5z�@�X���}�@`�c�aޜ@ �ԟ-K�@�AHD<�@�i8���BF������(@@�g�@ x�Z�j�@�/ con�@�R���Μ@ w�4�J�@���>�;�@�i8���BF`UUUU�(@����@ ���[�@����^�@ �/;��@ ��J�@ j��;�@�i8���BF     )@@O~�W��@@x1��L�@ �QbrO�@` �貯�@�%�*J�@@Y�I;�@�i8���BF�����*)@ p� ��@��y2x=�@ ����?�@ �]�0��@��Y��I�@�(4��:�@�i8���BFaUUUUU)@��;�`י@����W.�@�d~��0�@�򘏳��@�}��I�@�dʢ:�@�i8���BF    �)@���U�Ǚ@����<�@��Bl%!�@@��;��@ ��(I�@�MfmN:�@�i8���BF������)@��n���@���	'�@�t���@ ����q�@��"�H�@��j*�9�@�i8���BFbUUUU�)@@�����@���2�@��ºd�@@�4^b�@���zH�@�����9�@�i8���BF     *@@n����@ �`�@`Q���@`"�R�@��w#H�@ ��S9�@�i8���BF�����**@���a��@`����@ �u���@�ꦾ�C�@�s�v�G�@`χ 9�@�i8���BFcUUUUU*@@��{�@@U/�	Ԛ@��qԗ@��2?4�@ ��@tG�@�����8�@�i8���BF    �*@`�U�k�@���Ś@`k �*ŗ@����$�@�8�G�@@L��V8�@�i8���BF������*@��v\�@�(W���@`�֦굗@ �\^��@�H��F�@��K�8�@�i8���BFdUUUU�*@�ȏ4M�@��"-��@`�u尦�@�ډR�@`I}jF�@����7�@�i8���BF     +@@�_�=�@ �ЎD��@ =��}��@�*xI��@ ��F�@�N4`7�@�i8���BF�����*+@ KIi�.�@@���a��@`v�^Q��@ <ދ��@ �Y%�E�@���7�@�i8���BFeUUUUU+@ M����@����z�@ S�*y�@���؛@`@piE�@P �b�6�@�i8���BF    �+@�/�h�@@-�w�k�@�eӾ	j�@�$��tɛ@��_@E�@ #�ml6�@�i8���BF������+@@JC�D�@@�k��\�@�w���Z�@�YצK��@��6��D�@��L6�@�i8���BFfUUUU�+@@�'�@@��NN�@����K�@�~��)��@`H�mfD�@�?[$�5�@�i8���BF     ,@@��c�@�x�I?�@ ��<�@��(���@`���D�@P�)�~5�@�i8���BF�����*,@�KZ��Ә@�H��0�@����-�@�5ܙ���@��xȿC�@0U�15�@�i8���BFgUUUUU,@��^��Ę@`�	��!�@�о���@�ы�}�@���kC�@�U�=�4�@�i8���BF    �,@`���쵘@ �y5�@�	�$��@�����n�@� �6C�@3��4�@�i8���BF������,@`//!�@@F=�g�@�/��� �@���u�_�@ ���B�@@m��A4�@�i8���BFhUUUU�,@@^�@�r:���@@
-���@@�F��P�@ ���jB�@0dAd�3�@�i8���BF     -@�����@@8 ��@ ���@�'���A�@@���B�@`��]�3�@�i8���BF�����*-@����z�@�(��wؙ@�Ԗ@�3Z��2�@`��Y�A�@�L�Y3�@�i8���BFiUUUUU-@` fa(k�@��F��ə@`/Ŗ@ z�E$�@`9�DoA�@��)3�@�i8���BF    �-@@"��E\�@`5QqH��@ ��BU��@��� �@ ��A�@�wf�2�@�i8���BF������-@ �H�hM�@`�P����@ E����@ A�r>�@@�M��@�@�po2�@�i8���BFjUUUU�-@��>��>�@�S.��@�謲��@@���b��@���p@�@�m�Y"2�@�i8���BF     .@���o�/�@ ��.���@��4�ꉖ@��َ�@@��#@�@@c���1�@�i8���BF�����*.@ �k� �@��$�)��@`7){�@��(9�ٚ@�/��?�@p��*�1�@�i8���BFkUUUUU.@�쥥/�@��|,�r�@@�Dml�@��T��ʚ@ ��Sx?�@@QF�A1�@�i8���BF    �.@ ���o�@���~;d�@@hTh�]�@��#4��@���$?�@9��0�@�i8���BF������.@�8�����@�7m��U�@ �m�O�@��Zt��@�wh��>�@ Hb�0�@�i8���BFlUUUU�.@@�� �@`�b3aG�@@��iX@�@�9Ֆ���@���z>�@��x4[0�@�i8���BF     /@ 1��Qח@`W"��8�@ H�B�1�@@�R���@���w&>�@P�I�0�@�i8���BFª���*/@�G���ȗ@�.C(�*�@@�3#�@`YQL[��@�7���=�@ y���/�@�i8���BFmUUUUU/@������@�P�A�@`���w�@��&�r�@�T���=�@�B�|/�@�i8���BF    �/@�a��f��@�6�E��@ �q���@�n�td�@���,=�@��1/�@�i8���BFê����/@���lΜ�@�}�؛��@@rR��@�م�sU�@�����<�@��=U�.�@�i8���BFnUUUU�/@�8�o;��@`xv�P�@�]��@@��F�@��<�@�����.�@�i8���BF     0@@_��@@�?�
�@ �x�Cڕ@`��K8�@ ҆1<�@�贔R.�@�i8���BFaUUUU0@@�U�&q�@ �%.�Ԙ@�V���˕@�t߼�)�@��M��;�@�*&,.�@�i8���BF�����*0@`7��b�@ i��Ƙ@��?M��@�I�.=�@��� �;�@p���-�@�i8���BF    @0@ δq(T�@��2�X��@@i[�ٮ�@@I����@�:��:;�@ n`y-�@�i8���BF`UUUUU0@ �l��E�@ Q��'��@��Uk��@��{@��@�����:�@�<��.-�@�i8���BF�����j0@����?7�@�JFL���@ ���@�
b���@�(W�:�@�D�$�,�@�i8���BF
    �0@��:��(�@���Ӎ�@��?x���@@�5rY�@�d%?:�@�d�,�@�i8���BF_UUUU�0@�mRm�@����@����@u�@�����ҙ@ ��9�@�f�;V,�@�i8���BF������0@���W�@@-��q�@`R���f�@@�ę@����9�@&,�@�i8���BF	    �0@��aҰ��@�o9}c�@ ���X�@`'s�+��@ �\ H9�@@���+�@�i8���BF^UUUU�0@ iY�Z�@�*u&jU�@ �)HJ�@ �`VЧ�@�B?
�8�@ q^�}+�@�i8���BF������0@�/�	�@���[G�@@����;�@�΃�z��@�R�R�8�@���5+�@�i8���BF     1@ ��V�Җ@�5��R9�@@��˼-�@�?o�+��@�}NN8�@@����*�@�i8���BF]UUUU1@��}xĖ@ �}(O+�@`��!��@��wr�|�@�t�/�7�@�#N�*�@�i8���BF�����*1@@��:8��@`�F�P�@ �t(I�@ �AϠn�@�'܋�7�@�$O}f*�@�i8���BF    @1@�^+i���@��oW�@���3�@ �VRb`�@@��Z7�@@�2 *�@�i8���BF\UUUUU1@ !+�Ǚ�@ �(b�@�P�����@����'R�@ ��{7�@���)�@�i8���BF�����j1@ *�n���@�$K�q�@����@`���C�@�'�γ6�@ ����)�@�i8���BF    �1@�Bl}�@`񤁆�@@Є��ؔ@ � S�5�@`y,a6�@�]+�K)�@�i8���BF[UUUU�1@�H�rFo�@@��-�ח@`,�h�ʔ@ �Y@�'�@�T�6�@�5�)�@�i8���BF������1@�KD&a�@���ɗ@���i��@@-y�u�@ Ͼb�5�@�%L��(�@�i8���BF    �1@����
S�@�"T�⻗@ W1bW��@��m�V�@ �a}l5�@P*v�~(�@�i8���BFZUUUU�1@�!�D�@@��
��@ g�I��@�J�	<��@��ہ5�@ ���8(�@�i8���BF������1@�%
g�6�@��s�7��@�z�@��@ aC&�@@8�_�4�@�*~�'�@�i8���BF     2@ 2(��(�@�6ߕi��@�u�=��@@\K��@�_kt4�@p��'�@�i8���BFYUUUU2@������@`CX����@�u�w@v�@�}�9Ә@��$4�@ 5�n'�@�i8���BF�����*2@����@����v�@`���Hh�@�xjfŘ@��U�3�@`�*k,'�@�i8���BF    @2@@z����@��N�i�@�nYVZ�@`0����@�qă3�@@m���&�@�i8���BFXUUUUU2@ !���@ ��c[�@`��WhL�@ �����@�W��13�@��~E�&�@�i8���BF�����j2@`��W��@@+��M�@ ���~>�@`}k��@���2�@pbm�`&�@�i8���BF    �2@`��+Օ@�5È�?�@@䭚0�@  �*��@ ؠ}�2�@`�X�&�@�i8���BFWUUUU�2@�*Ǖ@�,��N2�@@If�"�@ ��@�@���y;2�@�,�D�%�@�i8���BF������2@�YWi:��@`�#V�$�@@n����@`�Dc[q�@�)�4�1�@�F3c�%�@�i8���BF    �2@ ��]��@ �z�@�.%��@@E�P{c�@@Z�s�1�@���Y%�@�i8���BFVUUUU�2@��Lb���@�|A*f	�@�0U\?��@���,�U�@�~��H1�@ @��%�@�i8���BF������2@�}$ⳏ�@`�S���@@�~�t�@�"���G�@���-�0�@�Z�.�$�@�i8���BF      3@`$j恕@`D�#7�@ ��ݓ@`� ��9�@ �٠�0�@p����$�@�i8���BFUUUUU3@ � t�@@��ۦ��@�cQO�ϓ@ eG�*,�@ �ӱT0�@�Y�S$�@�i8���BF�����*3@�b�[f�@��D�Ӗ@�2Z(5@ G��e�@`+��0�@@xs8$�@�i8���BF�����?3@ �sP�X�@ �8�Ŗ@�	0���@ g+,��@`Oqm�/�@�����#�@�i8���BFTUUUUU3@�a��J�@@���@�HyϦ�@@?�/��@ �|�e/�@P��ݔ#�@�i8���BF�����j3@`�0=�@ 4�N���@ lQ<#��@�lX/��@�bJ�/�@��WNS#�@�i8���BF�����3@@+���/�@�Z����@`x�{��@���{�@��>��.�@ �#�@�i8���BFSUUUU�3@ ���!�@ ��L���@ ���}�@���4�ٗ@`�slq.�@����"�@�i8���BF������3@�?��2�@`�e7��@@�==p�@���O%̗@ >~�!.�@����"�@�i8���BF������3@@q0���@�-�t�@���|�b�@��{4���@`�G�-�@���W"�@�i8���BFRUUUU�3@@������@�Q�feg�@���xU�@��@�Ⱇ@ �Ŗ�-�@`�!"�@�i8���BF������3@`�4�a�@��|�Z�@ ���G�@@���G��@�c�0-�@�Tt<�!�@�i8���BF������3@��.;�ݔ@�x�L�@�:ND�9�@�e�뱕�@  �
�,�@����!�@�i8���BFQUUUU4@ ���CД@`,��K?�@ Q�v,�@�}ys"��@@��,�@ '��\!�@�i8���BF�����*4@��{��@�)��1�@�_+o��@ `�,�z�@ {�PA,�@�'�;!!�@�i8���BF�����?4@ �:��@�7&<�$�@��2�}�@`���m�@��b �+�@�mC� �@�i8���BFPUUUUU4@@fs���@ ��[�@@&��@�JNܓ_�@�i��+�@�]ç �@�i8���BF�����j4@�~4E��@`�8�
�@� ���@�[jnR�@����R+�@���=i �@�i8���BF�����4@��Lь�@������@�d��+�@�����D�@`�.�+�@ �KC+ �@�i8���BFOUUUU�4@�^Xb�@����@�96K�ے@�:�*7�@@����*�@�3X���@�i8���BF������4@ ��J�q�@`��Y�@ )VKbΒ@�-�~�)�@�A��b*�@@N���@�i8���BF������4@@�3.�d�@ vS�#Օ@��Z��@��uU�@��_b*�@s��x�@�i8���BFNUUUU�4@@U�2W�@ Ӑ�Ǖ@@��񬳒@ E�J��@����)�@pr�<�@�i8���BF������4@���Y�I�@`��ź�@�p�X��@ A�ؐ�@���xt)�@P(����@�i8���BF������4@��w�<�@��7���@ K;D	��@���,5��@��$)�@p-����@�i8���BFMUUUU5@@�I�-/�@�1Ӣv��@�"Bx���@�
&���@ m�F�(�@��%���@�i8���BF�����*5@�/�/�!�@�S��@�l?�r~�@ C^q�ٖ@@$�ń(�@��>N�@�i8���BF�����?5@ �i���@`2��@����,q�@����7̖@@��24(�@ �P��@�i8���BFLUUUUU5@�S�(N�@ [�y�@���l�c�@@/�羖@��h)�'�@�fPJ��@�i8���BF�����j5@@R����@`I{�k�@���V�@���>���@��R`�'�@ ^�ޓ�@�i8���BF�����5@�2���@@����^�@��kI�@�АRM��@ ���3'�@P}[�R�@�i8���BFKUUUU�5@@�	�ߓ@�EuK�Q�@ �R2<�@����@ .x�&�@@X���@�i8���BF������5@�n�O[ғ@ ����D�@��f��.�@ T�dÉ�@�wZ��&�@P�W��@�i8���BF������5@ �W)œ@�i�`�7�@�`4:�!�@�\ά�|�@��W/&�@0��_��@�i8���BFJUUUU�5@ �m7���@`�ڮ*�@`�	��@ EE�Ko�@��Vi�%�@@H�U�@�i8���BF������5@ ���Ѫ�@�G���@�J^�x�@ [��b�@`��j~%�@`���@�i8���BF������5@`?�g���@���.��@@�B�T��@�F7��T�@���$%�@�a����@�i8���BFIUUUU6@�������@��Q��@@�P)5�@��=	�G�@�5b>�$�@`KĔ�@�i8���BF�����*6@���Ro��@�Ϸ��@ ?F���@�<���:�@`�u$�@��rW�@�i8���BF�����?6@`���Wv�@��ٺ��@��8�ӑ@ ��lj-�@@�?�$�@����@�i8���BFHUUUUU6@� }�Di�@�4(��ܔ@�=q��ő@���L �@ �<��#�@pS6���@�i8���BF�����j6@ ���6\�@ ���ϔ@�C��縑@`�r�0�@���3o#�@Pw�I��@�i8���BF�����6@ j��,O�@�8x�Ô@�]��ޫ�@�9�@���#�@`��t]�@�i8���BFGUUUU�6@@[�&B�@�z � ��@ �Eiڞ�@ ~�#��@`�}�"�@��&��@�i8���BF������6@@^��%5�@`1��A��@�t��ڑ�@������@�a�d"�@@�C���@�i8���BF������6@ v)(�@���Tg��@�W�7���@@�.>�ޕ@���"�@�`����@�i8���BFFUUUU�6@�:��1�@�<�����@ *�(�w�@ �ݫ�ѕ@��
L�!�@����h�@�i8���BF������6@ �VF>�@ �F����@���/�j�@�`Ay�ĕ@�Q��]!�@ ���*�@�i8���BF������6@ "�PO�@��(�u�@��DI
^�@�)�@ ���!�@p< ���@�i8���BFEUUUU7@�̴�d��@���%i�@ R�� Q�@��6����@�	ԃ� �@ ��*��@�i8���BF�����*7@@�?�~�@ u��_\�@@�w�<D�@�P�z��@���U �@�`�mu�@�i8���BF�����?7@@e���ڒ@ P�ݝO�@`�߈]7�@�����@�V�.  �@0|�;�@�i8���BFDUUUUU7@�vB��͒@�=j�B�@ {_�*�@��@i5��@`�Lq��@pH)]�@�i8���BF�����j7@@|�����@����&6�@�{�s��@��KQw�@ <�ZS�@��Mw��@�i8���BF�����7@�Y����@�P-q)�@ Zt���@@!,�oj�@����@�����@�i8���BFCUUUU�7@�1_E��@���=��@��@ ��]�@�gy���@���L�@�i8���BF������7@�6�/z��@ 1HZ�@`�z!A��@�Ǫ��P�@��K�@�S��@�i8���BF������7@�~+����@��o�g�@��z!|�@@�<��C�@ �*���@�?����@�i8���BFBUUUU�7@��LU�@��*���@����ݐ@�lQ7�@�Ֆ���@p�pA��@�i8���BF������7@�C�3t�@��ٔ �@�*P]�А@�i�GR*�@@���H�@05F�e�@�i8���BF������7@�&zg�@ /�Âݓ@@��FĐ@`�K���@ �����@P�.�*�@�i8���BFAUUUU8@�����Z�@ R��Г@���@��ǔ��@���k��@P�����@�i8���BF�����*8@�%�N�@�-�Rē@�e�O㪐@ [A�@���YC�@P�Aĸ�@�i8���BF�����?8@`���gA�@ ��R���@@�=�8��@@�G�V��@ ����@�+��@�i8���BF@UUUUU8@`�4�@@�W�3��@���Q���@�+��@ �Nv��@�)�bK�@�i8���BF�����j8@ ��(�@���z���@�i���@@����ݔ@�a�E�@P{e'�@�i8���BF�����8@@8�}�@��ʫ$��@�,5�Sx�@  �Iє@�U�/��@�����@�i8���BF?UUUU�8@��w���@`-"���@@*?w�k�@�cZ��Ĕ@@tE��@�9���@�i8���BF������8@�<��K�@@�k*$y�@�k��#_�@��6v���@�@�@�Ŷ!i�@�i8���BF������8@�}����@@���l�@�87ʒR�@`QW�`��@�G���@��t3�@�i8���BF>UUUU�8@�Coy+�@��)�3`�@���nF�@�*Ȟ�@��`���@P�SK��@�i8���BF������8@��¡ܑ@@��[�S�@�-h$~9�@ ��2��@ ��A�@��r��@�i8���BF������8@ ��9Б@@��RG�@`��,�@`��B���@���I��@@����@�i8���BF=UUUU9@ %њÑ@���:�@ �Fy �@�"��y�@���Ȕ�@�L�{W�@�i8���BF�����*9@��a���@ &���.�@`����@`�h�l�@�6�y?�@`��"�@�i8���BF�����?9@��eΤ��@@�;�"�@`����@����`�@�����@@�}n��@�i8���BF<UUUUU9@��Bk0��@�"޼��@@�n�&��@�ь��S�@ �Ҙ�@����@�i8���BF�����j9@���\���@����c	�@��@Jݏ@�¬G�@ J�E�@�FK���@�i8���BF�����9@�7qT��@ x�a��@�>�tď@ 6\Z�:�@�R����@�ݔ�P�@�i8���BF;UUUU�9@ 9���x�@ وs��@@�P���@ �..�@ �虙�@`�=�@�i8���BF������9@�J=��l�@���h�@�'ߒ�@`w�׭!�@@�"C�@���6��@�i8���BF������9@@�5�(`�@��/ؒ@��Z z�@ 2��@�@�����@����@�i8���BF:UUUU�9@`���S�@�(��˒@�i�ia�@@B�+��@�R����@@�e�y�@�i8���BF������9@�� �tG�@�*�o���@���ѺH�@ X�r��@@b�M@�@��6D�@�i8���BF������9@�y�� ;�@`nLJ��@ �e0�@@;L��@`Ea���@ �3��@�i8���BF9UUUU:@@>��.�@ Wm���@ �r�@��`��@��I���@�ƭ���@�i8���BF�����*:@`U�"�@�Ú�К�@ ������@�/�]Yד@@3Wu:�@0�Ψ��@�i8���BF�����?:@ Ku=�@��ݙ��@��CN�@�E�i˓@��@���@���q�@�i8���BF8UUUUU:@�ǭ��	�@@6)g��@�����͎@��C㸾�@ ����@pI�A�@�i8���BF�����j:@ �0����@ ��n8v�@��E�O��@ �eCo��@�6	�?�@� ��@�i8���BF�����:@�d���@@,[]j�@@��%ܜ�@���r(��@ j�y��@�����@�i8���BF7UUUU�:@ OM�H�@ 1���]�@���o��@@
��䙓@`�-:��@��s��@�i8���BF������:@ Ӎِ@�$��Q�@ W]!l�@@�;B���@�_&RA�@�rx9w�@�i8���BF������:@�DQ�̐@`��|�E�@@4/��S�@� k��@@rS���@��Y�F�@�i8���BF6UUUU�:@� �����@ e�'�9�@ b�];�@�bT6u�@ �mZ��@�c�V�@�i8���BF������:@��Q���@ M&�l-�@ ݡ#�@��si�@ Ֆ�H�@Д����@�i8���BF������:@ B��s��@@�f�W!�@ ��^�
�@@�Z��\�@�T���@`J_���@�i8���BF5UUUU;@ ��U��@���'F�@ 7�˔�@����P�@ ��p��@�1NQ��@�i8���BF�����*;@ h�;��@`��(8	�@��.aڍ@��_�D�@��1�M�@P�:/U�@�i8���BF�����?;@��؎$��@�I��-��@ �؟6@ Z�Hd8�@�<p���@@�'�@�i8���BF4UUUUU;@@��Ix�@ c�'�@ ��g��@ $8~H,�@`���@ fT9��@�i8���BF�����j;@ S�1l�@`�:%�@@�ם���@ ;Ө0 �@��C}Z�@pS����@�i8���BF�����;@����_�@ ��K&ّ@ ���y�@��z�@@@{��@`�9��@�i8���BF3UUUU�;@ �O��S�@ H�*͑@@�$��a�@ /���@ c)���@ `sn�@�i8���BF������;@ �D_�G�@�4�G2��@ �+��I�@ u����@�u@6b�@ #�5?�@�i8���BF������;@����;�@ைo=��@ �Q��1�@@s����@@����@�B��@�i8���BF2UUUU�;@���/�@��NL��@�H��@`�q���@�����@��:q��@�i8���BF������;@���q$�@ ���^��@@3Bd�@��i��ג@@�w)n�@��p8��@�i8���BF������;@�����@�9��t��@�q/�@����˒@����@`�7��@�i8���BF1UUUU<@`����@`�C=���@@��dBҌ@` F��@��6��@���]�@�i8���BF�����*<@�Q��4 �@ o��y�@ 5�m��@@y�l���@`���w�@@��~0�@�i8���BF�����?<@@4\ƚ�@�C� �m�@��+Q���@ kD��@ �b&�@�,/�@�i8���BF0UUUUU<@@u?�Џ@`�v$�a�@ ��܊�@ �x��@�����@��A��@�i8���BF�����j<@@����@`���V�@���|!s�@ �s�1��@ >���@�����@�i8���BF�����<@ ;2P_��@�kN+BJ�@@�j�m[�@���7L��@�&̼7�@POu��@�i8���BF/UUUU�<@��G���@ xٟp>�@ ~&ܿC�@�W��hx�@ ��C�
�@��Z�@�i8���BF������<@ P��r�@���7�2�@@xT�,�@��Hv�l�@��0�
�@p��-�@�i8���BF������<@��w'hZ�@@F�#�&�@@^6ry�@ ?F��`�@�þ�B
�@P!���@�i8���BF.UUUU�<@�G�o�B�@@xp��@��ء���@�����T�@ ����	�@p����
�@�i8���BF������<@�;ʇ>+�@`(�K�@@��"T�@��4kI�@�ώ�	�@@��
�@�i8���BF������<@�lXP��@`�Q:��@���͋@�� 4=�@ �ħS	�@�E\��
�@�i8���BF-UUUU=@�̮�3��@�
�����@ ;SOL��@��hg1�@�_{�	�@��9\
�@�i8���BF�����*=@�����@�����@�Kv�Ҟ�@����%�@ tb\��@p�J�1
�@�i8���BF�����?=@ vw�E͎@�xF)]��@ aH�`��@`�"g��@��ha�@@в�
�@�i8���BF,UUUUU=@@qJ�ڵ�@�A\�Ԑ@ �ڗ�o�@ ���@ o�x�@`y���	�@�i8���BF�����j=@ J�w��@��3��Ȑ@�/��X�@�lK_�@@^)���@`ƒ�	�@�i8���BF�����=@�o�Q��@ ��N��@�q��=A�@��!����@`�m}v�@�jb'�	�@�i8���BF+UUUU�=@�R��o�@ ������@�R��)�@`&
��@�X�&�@��C<k	�@�i8���BF������=@@��yX�@�E0: ��@�ܩW��@��*?ߑ@`+%��@�G�A	�@�i8���BF������=@�ݠ�3A�@`L��]��@ 5�X��@��/M�ӑ@ ��Ʌ�@�Mc�	�@�i8���BF*UUUU�=@��Ů�)�@ ��g���@@�Q�@ 
V�Ǒ@@�X�6�@��%I��@�i8���BF�����=@���k��@���"��@��%�̊@���@��@ A����@@�p���@�i8���BF������=@ aF����@�L�c�w�@���_���@�7^מ��@�YG���@�]p��@�i8���BF)UUUU>@��X6e�@�<�k�@������@఻G���@ �N,K�@0q&��@�i8���BF~����*>@�+m�C͍@ H\"c`�@�/<)p��@ _u�b��@�w2��@�u��X�@�i8���BF�����?>@�&��)��@�р;�T�@���Vp�@�9�2ʍ�@ �P��@p)�N2�@�i8���BF(UUUUU>@�;����@�+��HI�@�
p�EY�@ �E�6��@���*^�@��*�@�i8���BF}����j>@@|��@`ey��=�@@�4�<B�@ mYo�v�@ ����@�.����@�i8���BF�����>@ �A�q�@ �Q�<2�@�Y��;+�@���Uk�@�����@�_S��@�i8���BF'UUUU�>@@1*�Z�@ ��C�&�@�B�&A�@@d�n�_�@ �5w�@��.¡�@�i8���BF|�����>@@��$C�@����<�@ �5L��@ �T�@��|(�@ *|�{�@�i8���BF������>@�^�',�@`.w���@ �3�]�@`yT��H�@@����@���V�@�i8���BF&UUUU�>@@�S@�@ ��hI�@�=:/wω@��-=�@�����@ ��^2�@�i8���BF{�����>@�Ò�_��@�0�R��@��W����@���[�1�@`��>�@�O��@�i8���BF������>@�����@ T׃�ڏ@ �=����@@�$&�@ }h��@ � ��@�i8���BF
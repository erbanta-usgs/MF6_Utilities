cont double  40                                                                                        H3-13-8                                       �?q�#ɇ�#@UUUUUU�?ͅ{�Da#@�������?��	�(J#@�������?k�J��#@TUUUUU�?-̯Z�Y$@�������?�>�Ko$@�������?�
i��#@SUUUUU�?P�]%@#@�������?����#@�������?�n�A�#@RUUUUU�?-�f��N$@�������?�����$@�������?>$�}k-$@������ @�kv$��#@TUUUUU@p ��9#@������@w�&�#@������@Օ���3$@UUUUUU@cNۮ�y$@      @���
$@������@F���j#@VUUUUU@.�m#@     @��#��a#@������@+<�R$@WUUUUU@�]���$@     @�3z8Z$@������@:�-�#@XUUUUU	@ 쐔r=#@     
@�*�i#@������
@5|��$@YUUUUU@+�R-"w$@     @�rN{�F$@������@-�ǜ#@ZUUUUU@��\l.#@     @5h�k9#@������@�V��)�#@[UUUUU@_/�?�$@     @ժ�&M{$@XUUUUU@�����#@������@l�(�O#@     @�����M#@WUUUUU@5�C���#@������@B��$�e$@     @�	��
e$@VUUUUU@�R����#@������@��Ȯ4/#@      @��[Yy#@UUUUUU@��z�9�#@������@=��c$@������@�*s�$@TUUUUU@�;�S$@������@���
Bp#@������@��bM�=#@SUUUUU@�B�ç#@������@f�7]F$@������@����v$@RUUUUU@Az�\$@������@��g��V#@������@\��+�#@QUUUUU@}+��z#@������@���p7$@������@+�g��$@PUUUUU@���hHG$@������@��z���#@������@�š��:#@OUUUUU@^`8�{#@������@�0(�)$@������@����z$@NUUUUU@Axτ<5$@������@�e&7�#@������@^{���#@MUUUUU@��;U�K#@������@(f>�L$@������@{x\��$@LUUUUU@���n$@������@��y�#@������@����E#@KUUUUU@N��EZ#@������@-O"4�#@������@�2�p$@JUUUUU@��,Y$@������@Xn�魹#@������@I��0"#@IUUUUU@���<�)#@������@���5l�#@������@�NѱKu$@�����* @���,c�$@OUUUUU @`���#@����� @Y���_#@������ @ѧ��D#@PUUUU� @�r�r��#@������ @�兝W$@�����*!@/H�	�p$@QUUUUU!@�T�R}�#@�����!@6����C#@������!@$�ÿ'#@RUUUU�!@�Y�̏�#@������!@P6��M$@�����*"@3A��a�$@SUUUUU"@�#��1$@�����"@1�r��#@������"@(;��A;#@TUUUU�"@.)�*�#@������"@�5!�2$@�����*#@�Szqu{$@UUUUUU#@�H��$!$@     �#@L/6,o#@������#@�/^�#@VUUUU�#@ف#��`#@     $@�*���$@�����*$@�o��!�$@WUUUUU$@Q����]$@    �$@:�}�A�#@������$@��u�?#@XUUUU�$@v�C�]i#@     %@`�k�$@�����*%@" LMx$@YUUUUU%@�*��.J$@    �%@��<�'�#@������%@bU<k�#@ZUUUU�%@עd�8#@     &@b'��n�#@�����*&@��`�6�$@[UUUUU&@&y��}$@    �&@m4����#@������&@�9!�hQ#@\UUUU�&@82�sL#@     '@��հo�#@�����*'@��ʸc$@]UUUUU'@TR�&0e$@    �'@��,W�#@������'@���Q/#@^UUUU�'@�Ji\#@	     (@�h�j��#@�����*(@j&�[ _$@_UUUUU(@O����$@
    �(@Ą�}�$@������(@q	%A�o#@`UUUU�(@�}nQ�:#@     )@�C�DV�#@�����*)@�\jjqA$@aUUUUU)@-$)�`t$@    �)@�wB$@������)@�x�l$@bUUUU�)@<_�%�#@     *@��J���#@�����**@��UIq$@cUUUUU*@�R~ż�$@    �*@=O�^$@������*@�v�>��#@dUUUU�*@��CB#@     +@!w|�?}#@�����*+@"�:�!$@eUUUUU+@����z$@    �+@�|�6$@������+@��"V�#@fUUUU�+@ �XG#@     ,@�غ(�F#@�����*,@�!��#@gUUUUU,@NsH���$@    �,@�V��l$@������,@�8�#@hUUUU�,@"�G��C#@     -@�r˷vU#@�����*-@����-�#@iUUUUU-@l7y^l$@    �-@p"�[W$@������-@�ǆ�0�#@jUUUU�-@�r&) #@     .@)��Ť$#@�����*.@pp�G��#@kUUUUU.@�/�2�o$@    �.@��ؠ�$@������.@֧�[C�#@lUUUU�.@P�,�^#@     /@H٬a@#@ª���*/@bx��#@mUUUUU/@���!R$@    �/@a�0n$@ê����/@�����#@nUUUU�/@�9|�B#@     0@��=��#@aUUUU0@o����#@�����*0@:�>�G$@    @0@�O�$@`UUUUU0@	��R�0$@�����j0@�T��#@
    �0@n��=M7#@_UUUU�0@(��#@������0@�����,$@	    �0@��)��w$@^UUUU�0@]���$@������0@{w��m#@     1@�w}?7#@]UUUU1@��kGZ#@�����*1@�42$@    @1@��Z��$@\UUUUU1@�7;	\$@�����j1@v1
��#@    �1@U�!@<#@[UUUU�1@�0ԋ�c#@������1@;%� $@    �1@C�vNks$@ZUUUU�1@4��'H$@������1@�E|�#@     2@����#@YUUUU2@β�2#@�����*2@�@vWJ�#@    @2@�Q��}$@XUUUUU2@�~���{$@�����j2@c`��#@    �2@Z��'�O#@WUUUU�2@T��H#@������2@���Df�#@    �2@7��K`$@VUUUU�2@���-�d$@������2@�@_��#@      3@D�N0#@UUUUU3@��[#@�����*3@I���#@�����?3@/4�& \$@TUUUUU3@�>o��$@�����j3@Mav�$@�����3@���q#@SUUUU�3@j<��9#@������3@�����#@������3@�H7P1?$@RUUUU�3@����t$@������3@�R�E�$@������3@��1<X#@QUUUU4@>34�#@�����*4@byx-q#@�����?4@a��~�.$@PUUUUU4@}ha���$@�����j4@.����H$@�����4@�[1Ԁ�#@OUUUU�4@0g�_8#@������4@6Ë�Bt#@������4@��`�$@NUUUU�4@���>w$@������4@�滿o6$@������4@��z9w�#@MUUUU5@c��ۯ#@�����*5@�+�D#@�����?5@�5CG�#@LUUUUU5@���	�$@�����j5@���\o$@�����5@�*ŸV�#@KUUUU�5@�����F#@������5@ps�h�U#@������5@�9���#@JUUUU�5@\�+L�m$@������5@�7���[$@������5@���%��#@IUUUU6@�1]�$#@�����*6@qI�A=&#@�����?6@N����#@HUUUUU6@ʺ�Dq$@�����j6@���[+�$@�����6@T�P�^$@GUUUU�6@��R}Gc#@������6@!�8�B#@������6@-��a�#@FUUUU�6@�H"��S$@������6@%_�1Gr$@������6@>���#@EUUUU7@?LƽG#@�����*7@�"�Qi#@�����?7@l��/�#@DUUUUU7@�%邍H$@�����j7@���$@�����7@���Ϲ6$@CUUUU�7@G1�#@������7@ ��ԙ:#@������7@;����#@BUUUU�7@�g�-$@������7@���V{$@������7@sV���%$@AUUUU8@,�ix�s#@�����*8@����#@�����?8@��.{*[#@@UUUUU8@�M���$@�����j8@n�eʃ�$@�����8@��:	�a$@?UUUU�8@���A1�#@������8@��BZ@#@������8@Z
�+e#@>UUUU�8@]�Э� $@������8@�H�'v$@������8@�g�yM$@=UUUU9@\�t�#@�����*9@���#@�����?9@� ��M4#@<UUUUU9@F<r���#@�����j9@�Tp�$@�����9@����F�$@;UUUU�9@� �\�$@������9@!�"6O�#@������9@�_�(��#@:UUUU�9@����-"$@������9@���P�$@������9@���4�$@9UUUU:@3�ʊ�#@�����*:@���A#@�����?:@� p!�"#@8UUUUU:@�P��#@�����j:@|y�b�`$@�����:@^5�
��$@7UUUU�:@cUB�!$@������:@����x#@������:@�t9K�=#@6UUUU�:@~H��#@������:@BW�A$@������:@w�8�y$@5UUUU;@�4�}$@�����*;@�k�TP^#@�����?;@z��m+#@4UUUUU;@rN��q#@�����j;@ �t�/$@�����;@�Vn���$@3UUUU�;@T`��N$@������;@i�����#@������;@��Q�;#@2UUUU�;@wN�y�u#@������;@��2~�$@������;@��r�ez$@1UUUU<@���<$@�����*<@����#@�����?<@�䴮#@0UUUUU<@s���E#@�����j<@�n��#@�����<@��+Д�$@/UUUU�<@4;N-Is$@������<@�}��	�#@������<@p)��.I#@.UUUU�<@ ��_�U#@������<@��7���#@������<@�g�sm$@-UUUU=@h��]$@�����*=@��^SW�#@�����?=@2��u&#@,UUUUU=@ݧ�%#@�����j=@L��Q��#@�����=@Q�e|vo$@+UUUU�=@��G9�$@������=@E�0<$@������=@�`?;e#@*UUUU�=@�8<��A#@�����=@�����#@������=@�'�%�Q$@)UUUU>@��H�s$@~����*>@������#@�����?>@A���I#@(UUUUU>@�Rf�#@}����j>@�qs�#@�����>@��.��E$@'UUUU�>@V+����$@|�����>@b��O9$@������>@(ͨ 1�#@&UUUU�>@�7jrq:#@{�����>@6�+g�#@������>@f
\+$@
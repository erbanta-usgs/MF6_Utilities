cont double  40                                                                                        FLOW_1-5-6_1-6-6                              �?�վx"�@UUUUUU�?�3+��
�@�������?>3,b�@�������?�y����@TUUUUU�?s����@�������?O�^$��@�������?J.�=�@SUUUUU�?bf7� �@�������?.����%�@�������?�S�&$+�@RUUUUU�?��(s�0�@�������?}��U�6�@�������?n�!;=�@������ @�,	�E�@TUUUUU@�x�EJM�@������@ x,�U�@������@#vt8�^�@UUUUUU@�⋤�g�@      @&v-��q�@������@y؞f{�@VUUUUU@l�#���@     @`R��2��@������@#�0��@WUUUUU@.��T��@     @5@�屋@������@%"��P��@XUUUUU	@��%�}̋@     
@Y	��kً@������
@��=,�@YUUUUU@��w9��@     @��0����@������@< 0/�
�@ZUUUUU@�*��w�@     @%���!�@������@�k;�6-�@[UUUUU@Y!><8�@     @t��yC�@XUUUUU@j�N�@������@��T7�X�@     @�%�c�@WUUUUU@[�`^bn�@������@�
O�x�@     @Ay2;��@VUUUUU@�TfAr��@������@�Z�҅��@      @xYM�u��@UUUUUU@x��C��@������@�>���@������@���Rv��@TUUUUU@ǔ�B�ǌ@������@z�kь@������@�B�?ڌ@SUUUUU@9��%>�@������@�=���@������@�Ҝ��@RUUUUU@��/�n��@������@l�����@������@[k�/;�@QUUUUU@!��n�@������@������@������@�+�s&�@PUUUUU@1�E��.�@������@���y6�@������@{Da�V>�@OUUUUU@YP��F�@������@!���M�@������@��2YU�@NUUUUU@L}���\�@������@�[��5d�@������@�k��~k�@MUUUUU@�ˡ�r�@������@��T�y�@������@4�Bpɀ�@LUUUUU@~��۲��@������@���=���@������@(]�h=��@KUUUUU@U�a�ޛ�@������@�ZqNh��@������@�E�ڨ�@JUUUUU@�',N6��@������@��=:z��@������@_�s���@IUUUUU@T��3���@������@�|,�Ǎ@������@�LW�͍@�����* @P
1qӍ@OUUUUU @�R�>+ٍ@����� @��9;�ލ@������ @��?CZ�@PUUUU� @�=����@������ @j@�D/�@�����*!@��x�@QUUUUU!@ۈ�����@�����!@��W����@������!@��(���@RUUUU�!@�o���@������!@��[���@�����*"@�=����@SUUUUU"@�f��@�����"@�+��@������"@$����@TUUUU�"@��EJ�@������"@�����@�����*#@�"d�h!�@UUUUUU#@h�2e�#�@     �#@jw&�@������#@sF��I(�@VUUUU�#@�\^*�@     $@ٟl/X,�@�����*$@o��7.�@WUUUUU$@��/�@    �$@I%j�1�@������$@�73�@XUUUU�$@A.��4�@     %@�Ų-6�@�����*%@G��H7�@YUUUUU%@�2p8�@    �%@s�e�}9�@������%@O�q:�@ZUUUU�%@�'YfJ;�@     &@%:�h
<�@�����*&@rț��:�@[UUUUU&@p�vR9�@    �&@i�G�7�@������&@�i��6�@\UUUU�&@�ǒ65�@     '@�=̋�3�@�����*'@��@�s2�@]UUUUU'@Ac�1�@    �'@	Γ�/�@������'@�v�0I.�@^UUUU�'@8	8��,�@	     (@O���{+�@�����*(@6�V7*�@_UUUUU(@g�(�@
    �(@O!�C'�@������(@E���%�@`UUUU�(@&�0m$�@     )@���� #�@�����*)@
_�p�!�@aUUUUU)@�}�% �@    �)@��["��@������)@�w�G�@bUUUU�)@/�q���@     *@8��[e�@�����**@4H�"��@cUUUUU*@tlGd��@    �*@6Eb��@������*@�-"��@dUUUU�*@S�
�!�@     +@2M����@�����*+@��2�@eUUUUU+@��eT��@    �+@��K2A�@������+@������@fUUUU�+@��LK
�@     ,@c����@�����*,@��<IQ�@gUUUUU,@�й���@    �,@�I�rU�@������,@X�1J��@hUUUU�,@����U�@     -@0�7[���@�����*-@�Z�"R��@iUUUUU-@6�k}���@    �-@HJL��@������-@�K���@jUUUU�-@���B��@     .@�����@�����*.@��4��@kUUUUU.@.�(5��@    �.@�nH6%�@������.@X\�j���@lUUUU�.@���t�@     /@a��Y��@ª���*/@[ׯw��@mUUUUU/@E�)o�@    �/@g��j��@ê����/@;���T�@nUUUU�/@��d(��@     0@#+�B6�@aUUUU0@4�����@�����*0@��b��@    @0@Þ�/�ߍ@`UUUUU0@��;�ݍ@�����j0@l��:^܍@
    �0@��i�ڍ@_UUUU�0@6�5ٍ@������0@�����׍@	    �0@�r>�	֍@^UUUU�0@��Msԍ@������0@�?+��ҍ@     1@�JCэ@]UUUU1@×H��ύ@�����*1@�І΍@    @1@`��Nu̍@\UUUUU1@�����ʍ@�����j1@M�?ɍ@    �1@qB�Z�Ǎ@[UUUU�1@�U��ƍ@������1@'9�fč@    �1@�d�@ZUUUU�1@���()��@������1@�_R���@     2@��hS轍@YUUUU2@�j\F��@�����*2@�	㣺�@    @2@i�8��@XUUUUU2@>�J>^��@�����j2@參����@    �2@;x���@WUUUU�2@�p��o��@������2@7��ɰ�@    �2@eM{�"��@VUUUU�2@��{��@������2@��'ԫ�@      3@��nD+��@UUUUU3@e3hc���@�����*3@`���֦�@�����?3@II4,��@TUUUUU3@��N���@�����j3@�7)�ա�@�����3@=�d)��@SUUUU�3@���{��@������3@ʯk�͜�@������3@��eR��@RUUUU�3@�k�p��@������3@��!N���@������3@D�i��@QUUUU4@�Nc�_��@�����*4@��ʥ���@�����?4@���U���@PUUUUU4@j*7�H��@�����j4@|�����@�����4@Oh b⋍@OUUUU�4@1���-��@������4@	�C6x��@������4@>f_�@NUUUU�4@P�W��@������4@v��U��@������4@L2����@MUUUU5@�YK���@�����*5@�c |+~�@�����?5@�f�q|�@LUUUUU5@�z��z�@�����j5@�����x�@�����5@�>w@w�@KUUUU�5@O�a$�u�@������5@�U0��s�@������5@��5Y	r�@JUUUU�5@���Kp�@������5@�x8g�n�@������5@�Ɋ�l�@IUUUU6@<G�k�@�����*6@K�3�Mi�@�����?6@n�J��g�@HUUUUU6@�F$�e�@�����j6@�ُ	d�@�����6@�hGb�@GUUUU�6@l�Q�`�@������6@��L�^�@������6@Jy���\�@FUUUU�6@��_�6[�@������6@�w�qY�@������6@g@D�W�@EUUUU7@�z$��U�@�����*7@S�,T�@�����?7@�W�VR�@DUUUUU7@�~<ǍP�@�����j7@Rqj�N�@�����7@����L�@CUUUU�7@��I3K�@������7@P�ˀhI�@������7@$g�L�G�@BUUUU�7@dn���E�@������7@���6D�@������7@z�o,:B�@AUUUU8@��Lm@�@�����*8@�}&q�>�@�����?8@��d��<�@@UUUUU8@��`;�@�����j8@RR�M39�@�����8@�=d7�@?UUUU�8@�.�{�5�@������8@
���3�@������8@|�`�1�@>UUUU�8@5�� 0�@������8@� ��N.�@������8@�y5�|,�@=UUUU9@V����*�@�����*9@ ���(�@�����?9@0R�_'�@<UUUUU9@��w,%�@�����j9@x݋W#�@�����9@YL���!�@;UUUU�9@[
x���@������9@����@������9@�  �@:UUUU�9@B���(�@������9@p��Q�@������9@+�^�y�@9UUUU:@��ʩ��@�����*:@y[i��@�����?:@�:=C��@8UUUUU:@0ȣ�@�����j:@[A��8�@�����:@��6^�@7UUUU�:@�6-�	�@������:@S��'��@������:@}�d��@6UUUU�:@l����@������:@�7z��@������:@Y�0)2 �@5UUUU;@'?T��@�����*;@��u��@�����?;@c�K����@4UUUUU;@\^ֵ��@�����j;@�!����@�����;@*�n��@3UUUU�;@96b�@������;@eo��3�@������;@
�CR�@2UUUU�;@K)��o�@������;@�D�Ҍ�@������;@uPF��@1UUUU<@�a1��@�����*<@t�=k��@�����?<@cz����@0UUUUU<@D���@�����j<@��W4��@�����<@�k{Oތ@/UUUU�<@Ӄ��i܌@������<@�ǃڌ@������<@,A�،@.UUUU�<@�@౵֌@������<@���Ԍ@������<@�PX�Ҍ@-UUUU=@��^��Ќ@�����*=@��a1ό@�����?=@3�m-͌@,UUUUU=@MZ#Cˌ@�����j=@��XɌ@�����=@;�nǌ@+UUUU�=@�7���Ō@������=@	�VH�Ì@������=@�Ƌ���@*UUUU�=@�L�(ÿ�@�����=@z�?�ֽ�@������=@M�g�껌@)UUUU>@�Zp!���@~����*>@�!_��@�����?>@��b�#��@(UUUUU>@���5��@}����j>@L���F��@�����>@i�(=X��@'UUUU�>@�u��i��@|�����>@�Z��z��@������>@�*�x���@&UUUU�>@4�IO���@{�����>@Z᪪��@������>@���﹤�@
cont single                                                                                            L1DDN       L2DDN       fU8w�X��39��8��9X1B9�ME��N�9�0�9�u����::߀�9'�ɹ�o�:�p:�y���:�C,:�.����:\:�I_�xi;���:z���~�4;`�: |��A�a;�f�:<4ٺ�;��;X��lȫ;o�!;��#�/^�;PaE;�hG��N <�0p;�Wr��<ȑ;@ے��6=<ޚ�;����$�d<ח�;iGֻ�G�<M� <�����<��<�1����<'�;<�V:�&}�<��a<�c_�8	=@��<����..=̕�<�Ɵ�W�P=��<����Μy=�z�<`��v3�=�=���q�=H�*=P��2Q�=�M=:�<�]��=�Lv=]k^��>v�=7}��x�1>Ԑ�=�l���R>�.�=����w>���=��̽�Y�>?�>��%�><a8>ni����>�N]>�T��H�>�τ>͗'��?$f�>�8�i?	N�>��H���+?���>�V��A?��	?�]b�
�X?�U%?ńj�; p?.jF?��n���?Yn?z�n�y�?zߎ?�tj�K��?=t�?�nb�4�?[��?�4W��
�?~��?x|I�$��?�%@b�9�f��?